module full_test;
reg a;
reg b;
reg cin;
wire sum;
wire carry;
fulladder_task uut (.a(a), .b(b), .cin(cin), .sum(sum), .carry(carry));
initial
begin
$monitor($time,"a=%b b=%b cin=%b sum=%b carry=%b",a,b,cin,sum,carry);
a=0; b=0; cin=0;
#10 a=0; b=0; cin=1;
#10 a=0; b=1; cin=0;
#10 a=0; b=1; cin=1;
#10 a=1; b=0; cin=0;
#10 a=1; b=0; cin=1;
#10 a=1; b=1; cin=0;
#10 a=1; b=1; cin=1;
end
endmodule
